`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2019/06/24 09:26:51
// Design Name: 
// Module Name: csa
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module CSA_N_4#(parameter N = 222)(a,b,c,g,f);
input [N/3:0]a,b,c;
output [N/3:0]g,f;

assign g[0]=a[0]^b[0]^c[0];
assign g[1]=a[1]^b[1]^c[1];
assign g[2]=a[2]^b[2]^c[2];
assign g[3]=a[3]^b[3]^c[3];
assign g[4]=a[4]^b[4]^c[4];
assign g[5]=a[5]^b[5]^c[5];
assign g[6]=a[6]^b[6]^c[6];
assign g[7]=a[7]^b[7]^c[7];
assign g[8]=a[8]^b[8]^c[8];
assign g[9]=a[9]^b[9]^c[9];
assign g[10]=a[10]^b[10]^c[10];
assign g[11]=a[11]^b[11]^c[11];
assign g[12]=a[12]^b[12]^c[12];
assign g[13]=a[13]^b[13]^c[13];
assign g[14]=a[14]^b[14]^c[14];
assign g[15]=a[15]^b[15]^c[15];
assign g[16]=a[16]^b[16]^c[16];
assign g[17]=a[17]^b[17]^c[17];
assign g[18]=a[18]^b[18]^c[18];
assign g[19]=a[19]^b[19]^c[19];
assign g[20]=a[20]^b[20]^c[20];
assign g[21]=a[21]^b[21]^c[21];
assign g[22]=a[22]^b[22]^c[22];
assign g[23]=a[23]^b[23]^c[23];
assign g[24]=a[24]^b[24]^c[24];
assign g[25]=a[25]^b[25]^c[25];
assign g[26]=a[26]^b[26]^c[26];
assign g[27]=a[27]^b[27]^c[27];
assign g[28]=a[28]^b[28]^c[28];
assign g[29]=a[29]^b[29]^c[29];
assign g[30]=a[30]^b[30]^c[30];
assign g[31]=a[31]^b[31]^c[31];
assign g[32]=a[32]^b[32]^c[32];
assign g[33]=a[33]^b[33]^c[33];
assign g[34]=a[34]^b[34]^c[34];
assign g[35]=a[35]^b[35]^c[35];
assign g[36]=a[36]^b[36]^c[36];
assign g[37]=a[37]^b[37]^c[37];
assign g[38]=a[38]^b[38]^c[38];
assign g[39]=a[39]^b[39]^c[39];
assign g[40]=a[40]^b[40]^c[40];
assign g[41]=a[41]^b[41]^c[41];
assign g[42]=a[42]^b[42]^c[42];
assign g[43]=a[43]^b[43]^c[43];
assign g[44]=a[44]^b[44]^c[44];
assign g[45]=a[45]^b[45]^c[45];
assign g[46]=a[46]^b[46]^c[46];
assign g[47]=a[47]^b[47]^c[47];
assign g[48]=a[48]^b[48]^c[48];
assign g[49]=a[49]^b[49]^c[49];
assign g[50]=a[50]^b[50]^c[50];
assign g[51]=a[51]^b[51]^c[51];
assign g[52]=a[52]^b[52]^c[52];
assign g[53]=a[53]^b[53]^c[53];
assign g[54]=a[54]^b[54]^c[54];
assign g[55]=a[55]^b[55]^c[55];
assign g[56]=a[56]^b[56]^c[56];
assign g[57]=a[57]^b[57]^c[57];
assign g[58]=a[58]^b[58]^c[58];
assign g[59]=a[59]^b[59]^c[59];
assign g[60]=a[60]^b[60]^c[60];
assign g[61]=a[61]^b[61]^c[61];
assign g[62]=a[62]^b[62]^c[62];
assign g[63]=a[63]^b[63]^c[63];
assign g[64]=a[64]^b[64]^c[64];
assign g[65]=a[65]^b[65]^c[65];
assign g[66]=a[66]^b[66]^c[66];
assign g[67]=a[67]^b[67]^c[67];
assign g[68]=a[68]^b[68]^c[68];
assign g[69]=a[69]^b[69]^c[69];
assign g[70]=a[70]^b[70]^c[70];
assign g[71]=a[71]^b[71]^c[71];
assign g[72]=a[72]^b[72]^c[72];
assign g[73]=a[73]^b[73]^c[73];
assign g[74]=a[74]^b[74]^c[74];
    

assign  f[0]=(a[0]&b[0])|((a[0]^b[0])&c[0]);
assign  f[1]=(a[1]&b[1])|((a[1]^b[1])&c[1]);
assign  f[2]=(a[2]&b[2])|((a[2]^b[2])&c[2]);
assign  f[3]=(a[3]&b[3])|((a[3]^b[3])&c[3]);
assign  f[4]=(a[4]&b[4])|((a[4]^b[4])&c[4]);
assign  f[5]=(a[5]&b[5])|((a[5]^b[5])&c[5]);
assign  f[6]=(a[6]&b[6])|((a[6]^b[6])&c[6]);
assign  f[7]=(a[7]&b[7])|((a[7]^b[7])&c[7]);
assign  f[8]=(a[8]&b[8])|((a[8]^b[8])&c[8]);
assign  f[9]=(a[9]&b[9])|((a[9]^b[9])&c[9]);
assign  f[10]=(a[10]&b[10])|((a[10]^b[10])&c[10]);
assign  f[11]=(a[11]&b[11])|((a[11]^b[11])&c[11]);
assign  f[12]=(a[12]&b[12])|((a[12]^b[12])&c[12]);
assign  f[13]=(a[13]&b[13])|((a[13]^b[13])&c[13]);
assign  f[14]=(a[14]&b[14])|((a[14]^b[14])&c[14]);
assign  f[15]=(a[15]&b[15])|((a[15]^b[15])&c[15]);
assign  f[16]=(a[16]&b[16])|((a[16]^b[16])&c[16]);
assign  f[17]=(a[17]&b[17])|((a[17]^b[17])&c[17]);
assign  f[18]=(a[18]&b[18])|((a[18]^b[18])&c[18]);
assign  f[19]=(a[19]&b[19])|((a[19]^b[19])&c[19]);
assign  f[20]=(a[20]&b[20])|((a[20]^b[20])&c[20]);
assign  f[21]=(a[21]&b[21])|((a[21]^b[21])&c[21]);
assign  f[22]=(a[22]&b[22])|((a[22]^b[22])&c[22]);
assign  f[23]=(a[23]&b[23])|((a[23]^b[23])&c[23]);
assign  f[24]=(a[24]&b[24])|((a[24]^b[24])&c[24]);
assign  f[25]=(a[25]&b[25])|((a[25]^b[25])&c[25]);
assign  f[26]=(a[26]&b[26])|((a[26]^b[26])&c[26]);
assign  f[27]=(a[27]&b[27])|((a[27]^b[27])&c[27]);
assign  f[28]=(a[28]&b[28])|((a[28]^b[28])&c[28]);
assign  f[29]=(a[29]&b[29])|((a[29]^b[29])&c[29]);
assign  f[30]=(a[30]&b[30])|((a[30]^b[30])&c[30]);
assign  f[31]=(a[31]&b[31])|((a[31]^b[31])&c[31]);
assign  f[32]=(a[32]&b[32])|((a[32]^b[32])&c[32]);
assign  f[33]=(a[33]&b[33])|((a[33]^b[33])&c[33]);
assign  f[34]=(a[34]&b[34])|((a[34]^b[34])&c[34]);
assign  f[35]=(a[35]&b[35])|((a[35]^b[35])&c[35]);
assign  f[36]=(a[36]&b[36])|((a[36]^b[36])&c[36]);
assign  f[37]=(a[37]&b[37])|((a[37]^b[37])&c[37]);
assign  f[38]=(a[38]&b[38])|((a[38]^b[38])&c[38]);
assign  f[39]=(a[39]&b[39])|((a[39]^b[39])&c[39]);
assign  f[40]=(a[40]&b[40])|((a[40]^b[40])&c[40]);
assign  f[41]=(a[41]&b[41])|((a[41]^b[41])&c[41]);
assign  f[42]=(a[42]&b[42])|((a[42]^b[42])&c[42]);
assign  f[43]=(a[43]&b[43])|((a[43]^b[43])&c[43]);
assign  f[44]=(a[44]&b[44])|((a[44]^b[44])&c[44]);
assign  f[45]=(a[45]&b[45])|((a[45]^b[45])&c[45]);
assign  f[46]=(a[46]&b[46])|((a[46]^b[46])&c[46]);
assign  f[47]=(a[47]&b[47])|((a[47]^b[47])&c[47]);
assign  f[48]=(a[48]&b[48])|((a[48]^b[48])&c[48]);
assign  f[49]=(a[49]&b[49])|((a[49]^b[49])&c[49]);
assign  f[50]=(a[50]&b[50])|((a[50]^b[50])&c[50]);
assign  f[51]=(a[51]&b[51])|((a[51]^b[51])&c[51]);
assign  f[52]=(a[52]&b[52])|((a[52]^b[52])&c[52]);
assign  f[53]=(a[53]&b[53])|((a[53]^b[53])&c[53]);
assign  f[54]=(a[54]&b[54])|((a[54]^b[54])&c[54]);
assign  f[55]=(a[55]&b[55])|((a[55]^b[55])&c[55]);
assign  f[56]=(a[56]&b[56])|((a[56]^b[56])&c[56]);
assign  f[57]=(a[57]&b[57])|((a[57]^b[57])&c[57]);
assign  f[58]=(a[58]&b[58])|((a[58]^b[58])&c[58]);
assign  f[59]=(a[59]&b[59])|((a[59]^b[59])&c[59]);
assign  f[60]=(a[60]&b[60])|((a[60]^b[60])&c[60]);
assign  f[61]=(a[61]&b[61])|((a[61]^b[61])&c[61]);
assign  f[62]=(a[62]&b[62])|((a[62]^b[62])&c[62]);
assign  f[63]=(a[63]&b[63])|((a[63]^b[63])&c[63]);
assign  f[64]=(a[64]&b[64])|((a[64]^b[64])&c[64]);

assign  f[65]=(a[65]&b[65])|((a[65]^b[65])&c[65]);
assign  f[66]=(a[66]&b[66])|((a[66]^b[66])&c[66]);
assign  f[67]=(a[67]&b[67])|((a[67]^b[67])&c[67]);
assign  f[68]=(a[68]&b[68])|((a[68]^b[68])&c[68]);
assign  f[69]=(a[69]&b[69])|((a[69]^b[69])&c[69]);
assign  f[70]=(a[70]&b[70])|((a[70]^b[70])&c[70]);
assign  f[71]=(a[71]&b[71])|((a[71]^b[71])&c[71]);
assign  f[72]=(a[72]&b[72])|((a[72]^b[72])&c[72]);
assign  f[73]=(a[73]&b[73])|((a[73]^b[73])&c[73]);  

   assign  f[74]=(a[74]&b[74])|((a[74]^b[74])&c[74]);     
endmodule
